`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:55:13 04/26/2009 
// Design Name: 
// Module Name:    gpin_buf 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gpin_buf(
    input gpin0,
    input gpin1,
    input gpin2,
    input gpin3,
    input gpin4,
    input gpin5,
    input gpin6,
    input gpin7,
    input gpin8,
    input gpin9,
    input gpin10,
    input gpin11,
    input gpin12,
    input gpin13,
    input gpin14,
    input gpin15,
    input gpin16,
    input gpin17,
    input gpin18,
    input gpin19,
    input gpin20,
    input gpin21,
    input gpin22,
    input gpin23,
    input gpin24,
    input gpin25,
    input gpin26,
    input gpin27,
    input gpin28,
    input gpin29,
    input gpin30,
    input gpin31,
    output [31:0] gpin
    );

assign gpin[0] = gpin0;
assign gpin[1] = gpin1;
assign gpin[2] = gpin2;
assign gpin[3] = gpin3;
assign gpin[4] = gpin4;
assign gpin[5] = gpin5;
assign gpin[6] = gpin6;
assign gpin[7] = gpin7;
assign gpin[8] = gpin8;
assign gpin[9] = gpin9;
assign gpin[10] = gpin10;
assign gpin[11] = gpin11;
assign gpin[12] = gpin12;
assign gpin[13] = gpin13;
assign gpin[14] = gpin14;
assign gpin[15] = gpin15;
assign gpin[16] = gpin16;
assign gpin[17] = gpin17;
assign gpin[18] = gpin18;
assign gpin[19] = gpin19;
assign gpin[20] = gpin20;
assign gpin[21] = gpin21;
assign gpin[22] = gpin22;
assign gpin[23] = gpin23;
assign gpin[24] = gpin24;
assign gpin[25] = gpin25;
assign gpin[26] = gpin26;
assign gpin[27] = gpin27;
assign gpin[28] = gpin28;
assign gpin[29] = gpin29;
assign gpin[30] = gpin30;
assign gpin[31] = gpin31;

endmodule
