`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:10:51 04/26/2009 
// Design Name: 
// Module Name:    gpout_buf 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module gpout_buf(
    input [31:0] gpout,
    output gpout0,
    output gpout1,
    output gpout2,
    output gpout3,
    output gpout4,
    output gpout5,
    output gpout6,
    output gpout7,
    output gpout8,
    output gpout9,
    output gpout10,
    output gpout11,
    output gpout12,
    output gpout13,
    output gpout14,
    output gpout15,
    output gpout16,
    output gpout17,
    output gpout18,
    output gpout19,
    output gpout20,
    output gpout21,
    output gpout22,
    output gpout23,
    output gpout24,
    output gpout25,
    output gpout26,
    output gpout27,
    output gpout28,
    output gpout29,
    output gpout30,
    output gpout31
    );

assign gpout0 = gpout[0];
assign gpout1 = gpout[1];
assign gpout2 = gpout[2];
assign gpout3 = gpout[3];
assign gpout4 = gpout[4];
assign gpout5 = gpout[5];
assign gpout6 = gpout[6];
assign gpout7 = gpout[7];
assign gpout8 = gpout[8];
assign gpout9 = gpout[9];
assign gpout10 = gpout[10];
assign gpout11 = gpout[11];
assign gpout12 = gpout[12];
assign gpout13 = gpout[13];
assign gpout14 = gpout[14];
assign gpout15 = gpout[15];
assign gpout16 = gpout[16];
assign gpout17 = gpout[17];
assign gpout18 = gpout[18];
assign gpout19 = gpout[19];
assign gpout20 = gpout[20];
assign gpout21 = gpout[21];
assign gpout22 = gpout[22];
assign gpout23 = gpout[23];
assign gpout24 = gpout[24];
assign gpout25 = gpout[25];
assign gpout26 = gpout[26];
assign gpout27 = gpout[27];
assign gpout28 = gpout[28];
assign gpout29 = gpout[29];
assign gpout30 = gpout[30];
assign gpout31 = gpout[31];

endmodule
